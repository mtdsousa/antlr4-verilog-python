module hello();
    initial begin
        string s = "Hello";
        $display("%s", s);
    end
endmodule
