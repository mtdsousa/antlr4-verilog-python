module hello;
    string s = "Hello";
    initial begin
        $display("%s", s);
    end
endmodule
